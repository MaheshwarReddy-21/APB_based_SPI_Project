  
/********************************************************************************************

Copyright 2024 - Maven Silicon Softech Pvt Ltd.  
www.maven-silicon.com

All Rights Reserved.

This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd.
It is not to be shared with or used by any third parties who have not enrolled for our paid 
training courses or received any written authorization from Maven Silicon.

Filename                :       apb_defs.v   

module Name             :       ----

Description             :       Define files for APB based SPI Core testbench


*********************************************************************************************/

  `define APB_DATA_WIDTH 8
  `define SPI_REG_WIDTH 8
  `define APB_ADDR_WIDTH 3


